----------------------------------------------------------------------------------
-- Company:        
-- Engineer:       simon.burkhardt
-- 
-- Create Date:    2023-04-21
-- Design Name:    skid buffer testbench
-- Module Name:    tb_pattern_trig - bh
-- Project Name:   
-- Target Devices: 
-- Tool Versions:  GHDL 0.37
-- Description:    
-- 
-- Dependencies:   
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- this testbench acts as a streaming master, sending bursts of data
-- counting from 1-4, also asserting tlast on the 4th data packet

-- the testbench itself acts as a correct streaming master which keeps the data
-- until it is acknowledged by the DUT by asserting tready.

-- the data pattern can be influenced by the user in 2 ways
-- + Tx requests are generated by changing the pattern in p_stimuli_tready
--   the master will try to send data for as long as sim_valid_data = '1'
-- + Rx acknowledgements are generated by changing the pattern in p_stimuli_tready
--   the downstream slave after the DUT will signal ready-to-receive 
--   when sim_ready_data = '1'

-- simulate both with OPT_DATA_REG = True / False
entity tb_pattern_trig is
  generic
  (
    C_S_AXIS_TDATA_WIDTH  : integer := 512;
    C_COMPARE_DATA_WIDTH  : integer := 32
  );
end tb_pattern_trig;

architecture bh of tb_pattern_trig is
  -- DUT component declaration
  component pattern_detector is
    generic (
      C_S_AXIS_TDATA_WIDTH  : integer;
      C_COMPARE_DATA_WIDTH  : integer
    );
    port (
      AXIS_ACLK       : in  std_logic;
      AXIS_ARESETN    : in  std_logic;
      S_AXIS_TVALID   : in  std_logic;
      S_AXIS_TDATA    : in  std_logic_vector(C_S_AXIS_TDATA_WIDTH-1 downto 0);
      M_AXIS_TREADY   : in  std_logic;
      compare_pattern : in  std_logic_vector(C_COMPARE_DATA_WIDTH-1 downto 0);
      match_out       : out std_logic
    );
  end component;

  constant CLK_PERIOD: TIME := 5 ns;

  signal clk   : std_logic;
  signal rst_n : std_logic;


  signal o_s_axis_tvalid   : std_logic;
  signal o_s_axis_tdata    : std_logic_vector(C_S_AXIS_TDATA_WIDTH-1 downto 0);
  signal o_m_axis_tready   : std_logic;
  signal o_compare_pattern : std_logic_vector(C_COMPARE_DATA_WIDTH-1 downto 0);
  signal i_match_out       : std_logic;

  signal clk_count : std_logic_vector(7 downto 0) := (others => '0');
begin

  -- generate clk signal
  p_clk_gen : process
  begin
   clk <= '1';
   wait for (CLK_PERIOD / 2);
   clk <= '0';
   wait for (CLK_PERIOD / 2);
   clk_count <= std_logic_vector(unsigned(clk_count) + 1);
  end process;

  -- generate initial reset
  p_reset_gen : process
  begin 
    rst_n <= '0';
    wait until rising_edge(clk);
    wait for (CLK_PERIOD / 4);
    rst_n <= '1';
    wait;
  end process;

  -- accept and ack BRESP
  p_traffic_gen : process(clk)
  begin
    if rising_edge(clk) then
      if rst_n = '0' then
        o_s_axis_tdata <= (others => '0');
        o_m_axis_tready <= '1';
        o_s_axis_tvalid <= '0';
        o_compare_pattern <= x"deadbeef";
      else
        if unsigned(clk_count) = 5 then
          o_s_axis_tdata(511 downto 511-31) <= x"deadbeef";
          o_s_axis_tvalid <= '1';
        end if;
        if unsigned(clk_count) = 6 then
          o_s_axis_tdata <= (others => '0');
          o_s_axis_tvalid <= '0';
        end if;

        if unsigned(clk_count) = 12 then
          o_s_axis_tdata(511 downto 511-31) <= x"abababab";
          o_s_axis_tvalid <= '1';
        end if;
        if unsigned(clk_count) = 13 then
          o_s_axis_tdata <= (others => '0');
          o_s_axis_tvalid <= '0';
        end if;

        if unsigned(clk_count) = 17 then
          o_s_axis_tdata(511-32 downto 511-31-32) <= x"deadbeef";
          o_s_axis_tvalid <= '1';
        end if;
        if unsigned(clk_count) = 18 then
          o_s_axis_tdata <= (others => '0');
          o_s_axis_tvalid <= '0';
        end if;

      end if;
    end if;
  end process;

-- DUT instance and connections
  pattern_detector_inst : pattern_detector
    generic map (
      C_S_AXIS_TDATA_WIDTH  => C_S_AXIS_TDATA_WIDTH,
      C_COMPARE_DATA_WIDTH  => C_COMPARE_DATA_WIDTH
    )
    port map (
      AXIS_ACLK      => clk,
      AXIS_ARESETN   => rst_n,

      S_AXIS_TVALID   => o_s_axis_tvalid,
      S_AXIS_TDATA    => o_s_axis_tdata,
      M_AXIS_TREADY   => o_m_axis_tready,
      compare_pattern => o_compare_pattern,
      match_out       => i_match_out
    );

end bh;
